`include "main_tb.sv"
